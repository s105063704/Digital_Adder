module DBS();
  input clk;
  output reset;
  output data;
  
  always@() begin
    
  end
 
  
endmodule
