module DBS(good);
  input ;
  output ;
  output ;
  
  
endmodule
