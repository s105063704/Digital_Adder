module DBS();
  input ;
  output ;
  output ;
  
  
endmodule
