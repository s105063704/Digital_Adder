module DBS();
  input clk;
  output reset;
  output data_1;
  
  always@() begin
    
  end
 
  
endmodule
