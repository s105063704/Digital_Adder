module DBS();
  input clk;
  output reset;
  output data;
  
  
 
  
endmodule
