module DBS();

endmodule
