module DBS();
  input clk;
  output reset;
  output da;
  
  always@() begin
    
  end
 
  
endmodule
